
V1 7 0 dc 1V
V2 8 0 pwl (0 0V 1ns 1V)
V3 1 7 pwl (0 0V 1ns -1V)
R4 1 2 10
R5 8 9 10 

L1 2 3 192.94n
C1 3 4 100p
L2 9 10 192.94n
C3 10 6 100p
C4 10 4 100p

R3 0 5 10u
L3 5 4 192.94n

C2 3 6 100p
L0 7 6 192.94n

K01 L0 L1 0.155
K12 L1 L2 0.848
K23 L2 L3 0.155
K03 L0 L3 0.1
K02 L0 L2 0.155
K13 L1 L3 0.155


C12l 2 9 4.622p
C12r 3 10 4.622p




.tran 0.01ns 10ns 

.end

