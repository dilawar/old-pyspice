*Question 1_d: Decoupling

*Resistance
R1 1 2 50m
R2 0 5 50m

*Self Inductance
L1 2 3 1pH
L2 5 4 1pH

*Capacitance
C1 3 4 99nF
C2 6 4 1nF

Vdd 1 0 dc 1v
Ieq 3 6 PWL(0 0 50p 20 100p 0 1000p 0 1050p 20 1100p 0 2000p 0 2050p 20 2100p 0 3000p 0 3050p 20 3100p 0 4000p 0 4050p 20 4100p 0 5000p 0 5050p 20 5100p 0)
.ic v(3)=1
.tran 1ns 6ns uic

.control
	run
	plot  v(3)-v(4) 
.endc

.end 

