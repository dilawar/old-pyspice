*Question 3 , Assignment 2 

VDD 1 0 DC 1V

*Inductances Modelling

L11 1 2 195nH
L33 6 3 195nH
L44 0 4 195nH
L22 0 4 195nH
K13 L11 L33 0.152
K14 L11 L44 0.152
K12 L11 L22 0.0996
K34 L33 L44 0.837
K32 L33 L22 0.152
K42 L44 L22 0.152

*Capacitance Modelling

C13 2 3 104fF
C34 3 4 2.62pF
C42 4 4 104fF
C1 2 3 0.1n
C2 3 4 0.1n
R1 5 6 10

*Test voltage ramp
Vtest 5 0 PWL(0 0 1nS 1 50nS 1 1us 1 2us 1 3us) 


.tran 0.01ns 500ns uic
.control

run 
plot v(2) v(4)
.endc  
