*single ended signal

VDD a 0 DC 1V

R1 e f 10

L11 a b 195nH
L33 f c 195nH
L44 0 d 195nH
L22 0 d 195nH
K13 L11 L33 0.152
K14 L11 L44 0.152
K12 L11 L22 0.0993
K34 L33 L44 0.844
K32 L33 L22 0.152
K42 L44 L22 0.152

C1 b c 0.1n
C2 c d 0.1n
C13 b c 104.75fF
C34 c d 2.62pF
C42 d d 104.75fF

Vr e 0 PWL(0 0 1nS 1 50nS 1 1us 1 2us 1 3us) 

.tran 0.01ns 300ns uic
.control

run 
plot v(b) v(d)
.endc  
