*Question 3_b: Simple return path arrangement
*Resistance
R1 2 6 10

*Self Inductance
L1 1 3 193.7nH
L2 5 0 193.7nH
L3 6 4 193.7nH
L4 5 0 193.7nH

*Mutual Inductance
K13 L1 L3 0.1538
K14 L1 L4 0.1538
K12 L1 L2 0.1
K34 L3 L4 0.815
K32 L3 L2 0.1538
K42 L4 L2 0.1538

*Capacitance
C1 4 5 0.1nF
C2 3 4 0.1nF
C341 6 0 5.025pF
C342 4 5 5.025pF


Vdd 1 0 dc 1v
Vin 2 0 PWL(0 0 1ns 1 1us 1)
.tran 1ns 4ns uic

.control
	run
	plot v(3) v(5) 
.endc

.end 

