ques 3 part c


R1 9 10 10
R2 11 12 10

L1 3 4 0.248uH
L2 8 5 0.3882uH
L3 7 13 0.3882uH
L4 14 6 0.248uH

Ca 1 3 2.45pF
Cb 9 8 10.9pF
Cc 12 7 9.33pF
Cd 2 14 2.58pF

C1 4 5 0.1nF
C2 5 6 0.1nF
C3 4 13 0.1nF
C4 13 6 0.1nF


V1 1 0 1v
V3 1 10 pwl(0 0v 1ns 1v 2000ns 1v) 
V2 11 0 pwl(0 0v 1ns 1v 2000ns 1v)

.ic v(4)=1v v(6) = 0v
.tran 1ns 2000ns uic  
.end
