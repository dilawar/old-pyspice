Return path configuration

V1 1 0 DC 1.0V
V2 4 0 PWL(0 0 1ns 0 2ns 1 5ns 1 10ns 1) r = 5ns

R1 4 5 10
C1 2 3 0.1nf 
C2 3 6 0.1nf
.ic V(2) 0.01 v(3) 0.01
L11 1 2 0.194uH
L33 5 3 0.194uH
L44 0 6 0.194uH
L22 0 7 0.194uH
L31 3 2 29.83nH
L43 6 3 0.565uH
L21 7 2 19.502nH
L32 6 3 29.83nH
L41 6 2 29.83nH
L42 6 7 29.83nH

.tran 1n 50n uic



.end

