Q3.3 --- 09007021

.param Lset = 1e-10

Vin P Q dc 1V
V0 Q 0 dc 0v

L1 P R Lset
L2 Q S Lset

C1 A B 100n

R1 R A 5e-4
R2 S B 5e-4

.tran 1p 100ns uic
.plot v(a)-v(b)
.end
