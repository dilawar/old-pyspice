* Simulation for the peak ground-bounce and power-supply droop 
* at nodes R and S if a matched differential signaling
* arrangement is used in subsystems A and B

*Defining input voltage 
v1 1 0 1v

* Pulse r(t)with slope of 1 ns

vpulse1 1 3 pwl(0 0v 1ns 1v 50ns 1v)
vpulse2 6 0 pwl(0 0v 1ns 1v 50ns 1v)

* Defining self inductances
L11 1 2 193.348n
L33 4 5 193.348n

L44 7 8 193.348n 
L22 0 9 193.348n
*-----------------------------------------------------------
* Defining Mutual Inductances
K13 L11 L33 0.155
K14 L11 L44 0.155
K12 L11 L22 0.0999

K34 L33 L44 0.8483
K32 L33 L22 0.155

K42 L44 L22 0.155
*-----------------------------------------------------------
* Defining capacitances
C1 2 5 0.1n
C2 2 8 0.1n
C3 5 9 0.1n
C4 8 9 0.1n

*-----------------------------------------------------------
*Defining Resistances
R1 3 4 10
R2 6 7 10

------------------------------------------------------------
.tran 1ns 50ns 
 
* Control commands to run simulator, display the node status, and plot the specified results
.control

run

plot v(2)  
plot v(9)
set hcopydevtype=postscript
hardcopy differential_supplydroop.ps v(2) 
hardcopy differential_ground.ps v(9) 
.endc
* end Control commands

.end
