.TITLE ASSIGNMENT2 Q-3(b) PRASHANT SINGH 123070052
VDD	P	0 	DC	1
VRamp	1	V	PWL(0 0 1NS 1 2NS 1 5NS 1)
R1	1	U	10
CW101	P	0	0.88735PF
CW102	R	0	0.88735PF
CW341	U	V	4.62874PF
CW301	U	0	0.393615PF
CW401	V	0	0.51385PF
LW1	P	R	0.196731UH
LW2	Q	S	0.196731UH
LW3	U	W	0.196731UH
LW4	V	X	0.196731UH
KW3W4	LW3	LW4	0.8406
CW342	W	X	4.62874PF
CW302	W	0	0.393615PF
CW402	X	0	0.51385PF
CWX	W	X	0.1NF
CRW	R	W	0.1NF
CW201	Q	0	0.9206PF
CW202	S	0	0.9206PF
RGND	V	Q	0
RGND2	X	S	0
RGND3	Q	0	0
*use	tran	10ps	300ns in the command prompt
.end
	
