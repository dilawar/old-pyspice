*Que 3(c) modeling of the wires with for differnetial path arrangement



*************modelling the capacitances in the line******************************
C1 1 2 204.25ff
C2 4 5 204.25ff
C3 2 7 5.067pf	
C4 5 6 5.067pf
C5 7 0 204.25ff
C6 6 9 204.25ff

C7 4 5 100pf
C8 5 9 100ff
C9 4 10 100pf
C10 10 9 100pF
C11 2 0 204.25ff
C12 1 0 122.75ff
C13 6 9 204.75ff
C14 4 9 122.75ff
C15 7 1 204.25ff
C16 4 6 204.25ff

******************************** modelling the Self inductances********************
L1 1 4 192.315nH
L4 2 5 192.315nH
L3 7 6 192.315nH
L2 0 9 192.315nH

*****************************modelling the Mutual Inductances********************
K1 L1 L4 0.1544
K2 L4 L3 0.8534
K3 L3 L2 0.1544
K4 L2 L4 0.1544
K5 L3 L1 0.1544 

R1 2 3 10
R2 8 7 10
Vp 1 3 pwl(0 0v 1ns 1v 3ns 1v 70ns 1v)
Vq 8 0 pwl(0 0v 1ns 1v 3ns 1v 70ns 1v)

V1 1 0 1v

.tran 0.2ns 1us uic

.control

run

plot v(4) 
plot v(9)

plot v(4)-v(9)

.endc
.end
