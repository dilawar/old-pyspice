Assignment2 RollNo:113079011
*Matched differential signalling case

*Supply voltage
V1 	1	0 	dc 	1 
*Self inductances of the wires 			
L1	1	2	1.93564e-07		
L2	4	0	1.93564e-07		
L3	6	3	1.93564e-07		
L4	9	8	1.93564e-07	

*Coefficient of magnetic coupling between the wires
K12	L1	L2	0.0999819181 	
K34	L3	L4	0.84781261		
K14	L1	L4	0.153037238
K13	L1	L3	0.153120415
K23	L2	L3	0.153120415
K24	L2	L4	0.153037238


*Differential signals
V2	0	5	PWL(0 1 1n 0)
V3  1   11  PWL(0 0 1n 1)

*Differential signalling configuration
R1	5	9	10
R3  11  6   10
C1	2	8	0.1n
C2	2	3	0.1n
C3  3   4   0.1n
C4  8   4   0.1n

*Capacitance between Wire3 and 4(Split into two half value capacitors)
C5  6   9   4.80249e-12
C6  3   8   4.80249e-12

*Capacitance between Wire1 and 3(Split into two half value capacitors)
C7  1   6   2.04266e-13
C8  2   3   2.04266e-13

*Capacitance between Wire2 and 4(Split into two half value capacitors)
C9  9  0    2.04266e-13
C10  8   4   2.04266e-13

*Transient analysis duration
.TRAN 	0.1n	2000n


.end
*R2  7   0   10