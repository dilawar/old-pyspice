ques 1

v1 1 0 dc 1
r1 1 2 .5m
l1 2 3 0 
r2 0 4 .5m
l2 4 5 0
c1 3 5 99nf
c2 3 5 1nf


.tran .001ns 10ns uic
.end
