Question 3
*Circuit Description

Vdd P 0 dc 1V

*Inductances

L1  P R 1.9394e-7
L2  0 S 1.9394e-7
L3  U W 1.9394e-7
L4  V X 1.9394e-7

K12 L1 L2 0.1
K13 L1 L3 0.155
K14 L1 L4 0.155
K23 L2 L3 0.155
K24 L2 L4 0.155
K34 L3 L4 0.847


C1 R W 0.1e-9
C2 W X 0.1e-9

R1 1 U 10
R2 S X 0
R3 0 V 0

V1 1 V PWL(0 0 1ns 1 300ns 1)
.tran 1ns 300ns
.control
run
plot v(r) v(s)
.endc
.end
