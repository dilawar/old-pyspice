
Vdc 1 0 dc 1v
Vin 6 0 PWL(0 0 1ns 1V 10us 1V)  


C131 1 2 52.375f
C132 3 4 52.375f
C341 2 0 2.625p
C342 4 5 2.625p
C421 0 0 52.375f
C422 5 5 52.375f

C1 3 4 0.1n
C2 4 5 0.1n

R 3 2 10

L1 1 3 194nH
L2 0 5 194nH
L3 2 4 194nH
L4 0 5 194nH

K13 L1 L3 0.1543
K14 L1 L4 0.1504
K12 L1 L2 0.0358

K34 L3 L4 0.8434
K32 L3 L2 0.1543

K42 L4 L2 0.1543



.tran 1ns 2us uic

.control

run
plot v(3)
plot v(5)

.endc

.end 

