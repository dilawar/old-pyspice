assign23b

C13 1 3 200ff
*C15 1 5 200ff
*C10 1 0 120ff

C24 2 4 0.1nf
C26 2 6 0.1nf

C241 2 4 200ff
*C26 2 6 200ff
*C28 2 8 120ff

C35 3 5 5pf
*C30 3 0 200ff

C48 4 8 0.1nf

C46 4 6 5pf
*C481 4 8 200ff

C50 5 0 200ff
C68 6 8 200ff

C618 6 8 0.1nf

L12 1 2 193nH 
L34 3 4 193nH
L56 5 6 193nH
L08 0 8 193nH

K1234 L12 L34 0.154
*K1256 L12 L56 0.154
*K1208 L12 L08 0.100
K3456 L34 L56 0.854
*K3408 L34 L08 0.154
K5608 L56 L08 0.154

R1 7 3 10
R2 9 5 10


V10 1 0 1V

vina 1 7 PWL(0 0v 1ns 1v 5000.00ns 1v) 
vinb 9 0 PWL(0 0v 1ns 1v 5000.00ns 1v) 

.tran 0ns 5000ns

.control
run
plot v(8) v(2)
plot v(4) v(6)
.endc

.end