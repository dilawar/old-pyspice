DIFFERENTIAL SIGNAL CONFIGURATION

V1 1 0 dc 1.0V
V21 1 2 PWL(0 0 1ns 0 2ns 1 5ns 1 10ns 1) r=5ns
V22 5 0 PWL(0 0 1ns 0 2ns 1 5ns 1 10ns 1) r=5ns

L11 1 8  0.194uH  
L33 3 4  0.194uH  
L44 6 7  0.194uH
L22 0 9  0.194uH
L21 9 8  19.502nH
L32 9 4  29.83nH
L41 7 8  29.83nH  
L42 9 7  29.83nH
L43 7 4  0.565uH
L31 4 8  29.83nH
C3  9 4  0.1nf  
C1  4 8  0.1nf  
C4  9 7  0.1nf  
C2  7 8  0.1nf  
R1  2 3  10  
R2  5 6  10  

.ic v(8) 0.01 v(4) 0.01 v(7) 0.01

.tran 1n 50n uic

.end