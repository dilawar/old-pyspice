Vdd P 0 1V

L11 P R 195.8nH
L33 W U 195.8nH
L44 S 0 195.8nH
L22 S 0 195.8nH

K1 L11 L22 0.099101408
K2 L11 L33 0.152915828
K3 L11 L44 0.152831585
K4 L22 L33 0.152747342
K5 L22 L44 0.152830564
K6 L33 L44 0.835144132

C1 R W 0.1nF
C2 W S 0.1nF
R33 U M 10

VR M 0 pwl (0 0v 1ns 1v)
.tran 0.1ns 150ns uic
.control
run
plot v(R) v(S)
.endc
.end


