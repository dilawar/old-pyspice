

VDD 1 0 dc 1v
L1 1 8 .1942uH
L2 0 7 .1942uH
L3 3 5 .1942uH
L4 4 6 .1942uH 
R1 10 3 10
Vac 10 4 pwl(0ns 0v 1ns 1v 2ns 1v 3ns 1v 4ns 1v)
Vex 0 4 dc 0v
C1 5 8 0.1nf
C2 5 7 0.1nf
vex1 6 7 dc 0v



**mutual inductors

K1 L1 L2 .10008
K2 L3 L4 .80605
K3 L3 L1 .154682
K4 L4 L2 .154682
K5 L2 L3 .154682
K6 L1 L4 .154682

.ic v(8)=1v v(7)=0v v(5)=0v

.tran  0.1ns 1000ns uic
.end

 
