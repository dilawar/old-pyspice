* Simulation for the peak ground-bounce and power-supply droop at * nodes R and S if a return path arrangement is used in 
* subsystems A and B 

*Defining input voltage 
v1 1 0 1v

* Pulse r(t)with slope of 1 ns

vpulse 2 0 pwl(0 0v 1ns 1v 500ns 1v)

* Defining self inductances
L11 1 3 193.348n
L33 6 4 193.348n

L44 0 7 193.348n 
L22 0 5 193.348n
*-----------------------------------------------------------
* Defining Mutual Inductances
K13 L11 L33 0.155
K14 L11 L44 0.155
K12 L11 L22 0.0999

K34 L33 L44 0.8483
K32 L33 L22 0.155

K42 L44 L22 0.155
*-----------------------------------------------------------
* Defining capacitances
C1 3 4 0.1n
C2 4 7 0.1n
*-----------------------------------------------------------
*Defining Resistances
R1 2 6 10
R2 7 5 0.01
------------------------------------------------------------
.tran 1ns 500ns 
 
* Control commands to run simulator, display the node status, and plot the specified results
.control

run

plot v(3) v(5) 

set hcopydevtype=postscript
hardcopy returnpath.ps v(3) v(5)

.endc
* end Control commands

.end
