
*.MODEL custom_switch SW(VT=0.5v) 

Rdd 1 2 0.05
Rss 0 5 0.05

Cd 3 4 100nF 
 

L1 2 3 100nH 
L2 5 4 100nH 
v2 9 4 0v
V1 1 0 dc 1v
*I1 3 4 dc=0.5 pwl(0 0 0.95ns 0 1ns 10 1.05ns 0 1.95ns 0 2ns 10 2.0ns 0)
I1 3 9 dc=0.5 pulse(0 10 0 0.05ns 0.05ns 0.1ns 1ns)
.ic v(3) = 1v
.tran 1ns 10000ns uic
.end