Que 3(b) modeling of the wires with for return path arrangement

V1 1 0 1v

*************modelling the capacitances in the line******************************

C1 1 2 0.20425pf
C2 4 5 0.20425pf
C3 2 0 0.1925pf 
C4 5 7 0.1925pf
*C6 2 0 0.20425pf
*C7 1 0 0.122725pf
*C8 1 0 0.20425pf
*C9 7 5 0.20425pf
*C10 4 7 0.122725pf
*C11 4 7 0.20425pf
C12 4 5 0.1nf
C13 5 7 0.1nf

V2 6 7 0v


******************************** modelling the Self inductances********************

L1 1 4 0.192315uH
L4 2 5 0.192315uH
L3 6 0 0.192315uH
L2 7 0 0.192315uH

*****************************modelling the Mutual Inductances********************

K1 L1 L4 0.1544
K2 L1 L3 0.1544
K3 L4 L3 0.8534
K4 L4 L2 0.1544
K5 L3 L2 0.1544

R1 2 3 10
Vp 3 0 pwl(0 0v 1ns 1v 3ns 1v 70ns 1v)


.tran 0.2ns 10us uic

.control

run

plot v(4) 
plot v(3)
plot v(7)
plot v(4)-v(7)

.endc
.end
