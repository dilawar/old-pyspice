* Question 4b.

L1 1 2 1.933e-7
L2 4 3 1.933e-7
L3 0 6 1.933e-7
K L2 L3 1.6383e-7 

L4 0 6 1.933e-7
C1 3 6 8687ff
C2 2 3 0.1nf
C3 3 6 0.1nf
vin 1 0 1
vr1 5 0 pwl(0 0v 1ns 1v)


.tran .1ns 1000ns uic
.end


