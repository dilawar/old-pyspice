.include tsmc_spice_180nm.txt
R1 1 2 0.5m
C1 1 0 99n
C2 4 0 1n
L1 2 3 600u

v1 1 0 PWL(0 0 4.9n 0 5n 1 9.9n 1 10n 0);
v2 3 4 dc 0.0V
.tran 1n 10000n
.end